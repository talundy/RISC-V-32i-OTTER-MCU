`timescale 1ps / 1ns

module Stall(
	input clk,
	input rst,
	input rs1D,
	input rs2D,

	output logic stallF,
	output logic stallD,
	output logic flushE
	);





endmodule
